
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use std.textio.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity InstructionMemory is
    Port ( RST : in  STD_LOGIC;
           Address : in  STD_LOGIC_VECTOR (0 downto 31);
           instruction_out : out  STD_LOGIC_VECTOR (0 downto 31));
end InstructionMemory;

architecture Behavioral of InstructionMemory is
	type rom_type is array (63 downto 0) of std_logic_vector (31 downto 0);
	
	
	impure function InitRomFromFile (RomFileName : in string) return rom_type is
		FILE RomFile : text open read_mode is RomFileName;
		variable RomFileLine : line;
		variable temp_bv : bit_vector(31 downto 0);
		variable temp_mem : rom_type;
		begin
			for I in rom_type'range loop
				readline (RomFile, RomFileLine);
				read(RomFileLine, temp_bv);
				temp_mem(i) := to_stdlogicvector(temp_bv);
			end loop;
		return temp_mem;
	end function;
	
	signal instructions : rom_type := InitRomFromFile("testJMPL.data");
	
	
begin
	process(RST, Address,instructions)
	begin
			if(RST = '1')then
				instruction_out <= (others =>'0');
			else
				instruction_out <= instructions(conv_integer(Address(5 downto 0)));
			end if;
				
	end process;
end Behavioral;

